LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY tt_um_algorithmus_OSDungen IS
	PORT (
		clk : IN STD_LOGIC; -- 25 kHz
		reset: IN STD_LOGIC;
		p1_btn_left_in, p1_btn_right_in, p2_btn_left_in, p2_btn_right_in, start_btn_in : IN STD_LOGIC;
		leds_out : out STD_LOGIC_VECTOR(5 DOWNTO 0)
		  );
END tt_um_algorithmus_OSDungen;



ARCHITECTURE RTL OF tt_um_algorithmus_OSDungen IS

	COMPONENT RANDOM IS
		PORT (
			clk : IN STD_LOGIC;
			reset : IN STD_LOGIC;
			rnd_8bit_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) 
		);
	END COMPONENT;

    signal timer_counter: unsigned (16 downto 0);
    
    signal rnd_8bit : STD_LOGIC_VECTOR(7 DOWNTO 0); 
    
	TYPE t_state IS (s_reset, s_blinkOn1, s_blinkChange1, s_blinkOff1, s_blinkChange2, s_blinkOn2, s_blinkChange3,
	s_blinkOff2, s_blinkChange4, s_blinkOn3, s_blinkChange5, s_blinkOff3, s_waitRndInit, s_waitRnd, s_SetLeftLED,
	s_SetRightLED, s_P1Won, s_P2Won);
	SIGNAL state, next_state : t_state;
	
	signal timer_init_500msec, timer_decr, timer_init_rand: std_logic;
    
BEGIN

    I_RANDOM: component RANDOM
    port map (
      clk   => clk,
      reset => reset,
      rnd_8bit_out => rnd_8bit
    );


	-- Timer-Counter-Prozess (taktsynchroner Prozess)
	PROCESS (clk) -- (nur) Taktsignal in Sensitivitätsliste
	BEGIN
		IF rising_edge (clk) THEN
		    if (timer_init_500msec = '1') then
		         timer_counter <= "00011000100000000";
		    end if;

            if (timer_init_rand = '1') then
				timer_counter <= unsigned(rnd_8bit(2 downto 0) & "11000100000000");
			end if;
		        
		    if (timer_decr = '1') then
                timer_counter <= timer_counter - 1;
            end if;
		END IF;
	END PROCESS;

	-- Zustandsregister (taktsynchroner Prozess)
	PROCESS (clk) -- (nur) Taktsignal in Sensitivitätsliste
	BEGIN
		IF rising_edge (clk) THEN
		    IF (reset = '1') then
		        state <= s_reset;
		    ELSE
			    state <= next_state;
			END IF;
		END IF;
	END PROCESS;
	

	-- Prozess für die Uebergangs- und Ausgabefunktion
	PROCESS (state, p1_btn_left_in, p1_btn_right_in, p2_btn_left_in, p2_btn_right_in, start_btn_in, rnd_8bit, timer_counter) -- Zustand und alle Status-Signale in Sensitiviaetsliste 
	BEGIN
	
	    timer_init_500msec <= '0';
	    timer_init_rand <= '0';
	    timer_decr <= '0';
	    
	    leds_out <= (others => '0');
	    
	    next_state <= state;
	    
		CASE state IS
			WHEN s_reset =>
				IF start_btn_in = '1' THEN
					next_state <= s_blinkOn1;
				END IF;
				
				timer_init_500msec <= '1';			
				
			WHEN s_blinkOn1 =>
				leds_out <= (others => '1');
				
				if timer_counter = 0 then
					next_state <= s_blinkChange1;
				else
				    timer_decr <= '1';
				end if;
			
			WHEN s_blinkChange1 =>
				timer_init_500msec <= '1';
				next_state <= s_blinkOff1;
			
			WHEN s_blinkOff1 =>
				leds_out <= (others => '0');
				
				if timer_counter = 0 then
					next_state <= s_blinkChange2;
				else
				    timer_decr <= '1';
				end if;
			
			WHEN s_blinkChange2 =>
				timer_init_500msec <= '1';
				next_state <= s_blinkOn2;
			
			WHEN s_blinkOn2 =>
				leds_out <= (others => '1');
				
				if timer_counter = 0 then
					next_state <= s_blinkChange3;
				else
				    timer_decr <= '1';
				end if;
			
			WHEN s_blinkChange3 =>
				timer_init_500msec <= '1';
				next_state <= s_blinkOff2;
			
			WHEN s_blinkOff2 =>
				leds_out <= (others => '0');
				
				if timer_counter = 0 then
					next_state <= s_blinkChange4;
				else
				    timer_decr <= '1';
				end if;
			
			WHEN s_blinkChange4 =>
				timer_init_500msec <= '1';
				next_state <= s_blinkOn3;
			
			WHEN s_blinkOn3 =>
				leds_out <= (others => '1');
				
				if timer_counter = 0 then
					next_state <= s_blinkChange5;
				else
				    timer_decr <= '1';
				end if;
				
			WHEN s_blinkChange5 =>
				timer_init_500msec <= '1';
				next_state <= s_blinkOn3;
				
			WHEN s_blinkOff3 =>
				leds_out <= (others => '0');
				
				if timer_counter = 0 then
					next_state <= s_waitRndInit;
				else
				    timer_decr <= '1';
				end if;

			WHEN s_waitRndInit => 
			    timer_init_rand <= '1';
			    next_state <= s_waitRnd;
			
			WHEN s_waitRnd =>
			    timer_decr <= '1';
			    
				IF timer_counter = 0 THEN
					if rnd_8bit(7) = '1' then
						next_state <= s_SetLeftLED;
					else
						next_state <= s_SetRightLED;
					end if;
				ELSIF p1_btn_left_in = '1' or p1_btn_right_in = '1' then 
					next_state <= s_p2Won;
				ELSIF  p2_btn_left_in = '1' or p2_btn_right_in = '1' then 
					next_state <= s_p1Won;
				END IF;

			WHEN s_SetLeftLED =>
				leds_out(0) <= '1';
				if (p1_btn_left_in = '1' or p2_btn_right_in = '1') then
					next_state <= s_P1Won;
				elsif (p1_btn_right_in = '1' or p2_btn_left_in = '1') then
					next_state <= s_P2Won;
				end if;
					
			WHEN s_SetRightLED =>
				leds_out(1) <= '0';
				if (p1_btn_right_in = '1' or p2_btn_left_in = '1') then
					next_state <= s_P1Won;
				elsif (p1_btn_left_in = '1' or p2_btn_right_in = '1') then
					next_state <= s_P2Won;
				end if;

			WHEN s_P1Won =>
			    leds_out(3 downto 2) <= "11";
				timer_init_500msec <= '1';	
				
			    if start_btn_in = '1' then
					next_state <= s_blinkOn1;
				end if;

			WHEN s_P2Won =>
			    leds_out(5 downto 4) <= "11";
				timer_init_500msec <= '1';	
				
			    if start_btn_in = '1' then
					next_state <= s_blinkOn1;
				end if;
		END CASE;
	END PROCESS;
END RTL;
